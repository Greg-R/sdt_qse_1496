* 2nd Stage of the SDT Transmitter

.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/2N3904.LIB"
*.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/MMBT2222ALT1.LIB"

.subckt amplifier2 input output vsupply
* NPN BJT Collector Base Emitter
Q2 output 2 3 Q2n3904

C2 input 2 0.2u
Rconverge input 0 2.0Meg

R5  2 0 3300.0
R6  output 2 5600.0
R7  vsupply output 1200.0
R8  3 0    100.0
C4  3 0    0.390p

L1   vsupply 4      0.18u
R10  4       5      680.0
C3   5       output 0.1u


.ends amplifier2