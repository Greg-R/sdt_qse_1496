Simulate MC1496 based IQ Modulator
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_xmas_travel/MC1496_SPICE_MODEL.LIB"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_xmas_travel/MMBT2222ALT1.LIB"

.subckt dsbmodulator audioin rfin outplus outminus
.param loadrf = 1000 bullshit = 1000
Vsupply 15 0 DC 12.27 
* MC1496 VS+ GAIN2 GAIN3 VS- Bias VO+ NC VEE NC VO- NC VC- NC VC+
XGCELL    1    2 3 4 5 6 7 0 9 12 11 10 13 8 MC1496
* Output bias resistors
Rloadplusi   15  6 3000
Rloadminusi  15 12 3000
* Gain setting resistor
Rgain 2 3 1000
* Main bias control resistor
Rbias 15 5 10000
* Bias chain
R1 15  8 1300
R2  8 17  820
R3 17  0 1000
* Signal input bias
R4 17 1 1000
R5 17 4 1000
* Signal input blocking capacitor
C1i audioin 1 0.1u
* Signal bypass capacitors, for both RF and audio.
Caudiobypassi 4 0 100.0u ic=3.905v
Crfbypassi 8 0 100.0u ic=7.135v
* Carrier input bias
R6i 8 10 51
* RF input blocking capacitor
C2i rfin 10 0.1u

* Output emitter followers and blocking caps.
Qoutplusi  15 6 120 Qmmbt2222alt1g
Qoutminusi 15 12 121 Qmmbt2222alt1g
Rlplusi 120 0 1000 
Rlminusi 121 0 1000 
Coutplusi 120 outplus 0.1u
Coutminusi 121 outminus 0.1u

.ends dsbmodulator

xmodi 1 2 outplusi outminusi dsbmodulator
xmodq 3 4 outplusq outminusq dsbmodulator

.param audiolevel = 400.0m lolevel = 150.0m
.param rffreq = 7.0e6

Viaudio 1 0 sin(0 {audiolevel} 1000 0.1m 0 0)
Vilo    2 0 sin(0.0, {lolevel}, {rffreq}, 0.1m, 0 0)
Vqaudio 3 0 sin(0 {audiolevel} 1000 0.1m 0 90)
Vqlo    4 0 sin(0.0, {lolevel}, {rffreq}, 0.1m, 0, 90)

* Join the positive outputs together with small resistors.
Rplusi outplusi outplus 1.0
Rplusq outplusq outplus 1.0
*Rloadplus outputplus 0 loadrf

* Join the negative outputs together with small resistors.
Rminusi outminusi outminus 1.0
Rminusq outminusq outminus 1.0
*Rloadminus outputminus 0 loadrf

* A transformer on the outout.
Lprimary outplus outminus 1000u
Lsecondary output 0 70u
Ktrans Lprimary Lsecondary 1.0

* RF Load
Rload output 0 50.0

.control
set ngbehavior=ps

if i > 0
echo {$&i}
else
let i = 0
end

compose secondary values 100u 200u 400u 700u 1000u 1500u 2000u 2770u 4000u 6000u
let fundmag = vector(10)

*destroy all
save output

while i < 10
alter Lsecondary = secondary[i]
tran 10.0n 15.1m 10.1m uic
*setplot tran1
*plot output

*setplot tran1
*  Try Fourier analysis.
fourier 7.0Meg v(output)
let i = i + 1
*plot fourier{$&i}1[1] vs fourier{$&i}1[0]
let j = i - 1
let fundmag[{$&j}] = fourier{$&i}1[1][1]
end

plot fundmag vs secondary

*compose fundmag values fourier11[1][1] fourier21[1][1] fourier31[1][1]

*destroy all
*setplot tran1
*linearize output
*set specwindow = blackman 
*fft output
*plot db(output) xlimit 6.995e6 7.005e6  ylimit -100 0.0 ydelta 10.0
*plot db(output) ylimit -100.0 0.0 ydelta 10.0

.endc

.end
