* Simulation of a simple BJT cascode amplifier for HF.
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/MMBT2222ALT1.LIB"

.MODEL Q_JS04_N_1 NPN( IS=9.99F NF=1 NR=1 RE=2.51 RC=1 
+      RB=10 VAF=40 VAR=20 ISE=4.03P ISC=4.03P 
+      ISS=0 NE=1.78 NC=1.78 NS=1 BF=679 
+      BR=5 IKF=13.8M IKR=13.8M CJC=3.6P CJE=3.99P 
+      CJS=0 VJC=878M VJE=16.1 VJS=750M MJC=307M 
+      MJE=2.01 MJS=0 TF=531P TR=69N EG=1.11 
+      KF=0 AF=1 )
.END

Vsupply 12 0 DC 12.0V

Qce 1 2 3 Q_JS04_N_1
Qcb 4 5 1 Q_JS04_N_1

* Emitter resistor
Re 3 0 0.1
* Bias the base of the CE amp.
R1 12 2 10000.0
Rb 2  0  1539.0
* Bias the base of the CB amp.
R2 12 5  5000.0
Rcb 5 0  5000.0
* AC shunt the base to ground.
Cbase 5 0 10.0u

Rl 12 4   500.0

* Input and output blocking capacitors.
Cin input   2 1.0u
Cout output 4 1.0u
* Load resistors
Rin input   0 1.0Meg
Rout output 0 1000.0

Vin input 0 DC 0 AC 1

.control
set ngbehavior=ps

ac dec 10 1000 100.0e6

plot db(v(output))
plot db(v(1))

.endc

.end


