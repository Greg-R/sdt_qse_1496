* MC1496 based DSB Modulator
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/MC1496_SPICE_MODEL.LIB"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/MMBT2222ALT1.LIB"

.subckt dsbmodulator audioin rfin 18 19

Vsupply 15 0 DC 12.27
Vhigh  22 0 DC 24.0
* MC1496 VS+ GAIN2 GAIN3 VS- Bias VO+ NC VEE NC VO- NC VC- NC VC+
XGCELL    1    2     3    4   5    6  7   0  9  12  11 10  13  8  MC1496
* Output bias resistors
*Rloadplusi   15  6 1000
*Rloadminusi  15 12 1000
* Gain setting resistor
Rgain 2 3 500
* Main bias control resistor
Rbias 15 5 10000
* Bias chain
R1 15  8 1300
R2  8 17  820
R3 17  0 1000
* Signal input bias
R4 17 1 100
R5 17 4 100
* Signal input blocking capacitor
C1i audioin 1 1.0u ic=-3.918
* Signal bypass capacitors, for both RF and audio.
Caudiobypassi 4 0 10.0u ic=3.918v
Crfbypassi 8 0 10.0u ic=7.20v
* Carrier input bias
R6i 8 10 51
* RF input blocking capacitor
C2i rfin 10 0.1u

*  Temporary output blocking capacitors
*Coutplusi  18 outplus 0.1u
*Coutminusi 19 outminus 0.1u
*Routplusi  outplus  0 1.0Meg
*Routminusi outminus 0 1.0Meg

* Output cascodes and blocking caps.
Qoutplus   18 20  6 Qmmbt2222alt1g
Qoutminus  19 21 12 Qmmbt2222alt1g
Rlplusi    22 18 1000.0
Rlminusi   22 19 1000.0
Rbias1     15 20 400.0
Rbias2     20  0 1000.0
Rbias3     15 21 400.0
Rbias4     21  0 1000.0
Cbypassplus  20 0 0.2u
Cbypassminus 21 0 0.2u
*Coutminusi 121 outminus 0.1u
*Routplusi  outplus 0 1.0Meg
*Routminusi outminus 0  1.0Meg

* Output emitter followers and blocking caps.
*Qoutplusi  15 6 120 Qmmbt2222alt1g
*Qoutminusi 15 12 121 Qmmbt2222alt1g
*Rlplusi    120 0 1000 
*Rlminusi   121 0 1000 
*Coutplusi  120 outplus 0.1u
*Coutminusi 121 outminus 0.1u
*Routplusi  outplus 0 1.0Meg
*Routminusi outminus 0  1.0Meg

.ends dsbmodulator
