* 2nd Stage of the SDT Transmitter

* Include the sub-circuit.
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_original/simulation_second_stage/second_stage_amp_subckt.cir"

* Needs a 15 volt power source:
Vsupply vsupply 0 15V

* Connect the output of the first stage to the base of the second stage.
Xfirststage input output vsupply amplifier2

.param rflevel = 150.0m
.param rffreq = 7.0e6

* Input source
Vin input 0 sin(0 {rflevel} {rffreq} 0.1m 0 0)

* Input source
*Vin 1 0 dc 0 ac 1.0 portnum 1 z0 50.0
* Output source
*Vout 2 0 dc 0 ac 1.0 portnum 2 z0 50.0

.control
set ngbehavior=ps
*save input output
*op
*ac dec 10 1.0Meg 100.0Meg
*sp dec 10 1.0Meg 100.0Meg

tran 2n 1.1m 1.099m

plot v(output)
plot v(input)
.endc

.end