* 2nd Stage of the SDT Transmitter

* Include the sub-circuit.
*.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_2N3904_amp/amplifier_2n3904.cir"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_2N3904_amp/2N3904.LIB"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_xmas_travel/MMBT2222ALT1.LIB"
* Include the sub-circuit.
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_2N3904_amp/amplifier_2n3904.cir"

* Needs a 15 volt power source:
Vsupply 15 0 15V

* Connect the output of the first stage to the base of the second stage.
Xfirststage firstin secondin 15 amplifier

Rloadfirst secondin 14 50.0
Cblock 14 0 0.1u

* Instantiate a transistor C B E
Q2 1 secondin 3 Qmmbt2222alt1g

R7 15 1 1200
R6  1 secondin 5600
R5  secondin 0 3300
R8  3 0  200
Co  1 output 0.1u
Rloadsecond output 0 5000

.param rflevel = 150.0m
.param rffreq = 7.0e6

* Input source
Vin firstin 0 sin(0 {rflevel} {rffreq} 0.1m 0 0)

* Input source
*Vin 1 0 dc 0 ac 1.0 portnum 1 z0 50.0
* Output source
*Vout 2 0 dc 0 ac 1.0 portnum 2 z0 50.0

.control
set ngbehavior=ps
save secondin output
*op
*ac dec 10 1.0Meg 100.0Meg
*sp dec 10 1.0Meg 100.0Meg

tran 10n 1.1m 1.0m

plot v(output)
plot v(secondin)
.endc

.end