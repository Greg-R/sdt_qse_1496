Simulate MC1496 based IQ Modulator
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_iq_modulator/dsbmod_subckt.cir"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/feedback_amp_subckt.cir"

Vsupply 15 0 DC 12.27

xmodi 1 2 30 31 15 dsbmodulator
xmodq 3 4 30 31 15 dsbmodulator

* DSB modulator output bias resistors
Rbiasi 15 30 500.0
Rbiasq 15 31 500.0

.param audiolevel = 200.0m lolevel = 100.0m
.param rffreq = 28.0e6

Viaudio 1 0 sin(0 {audiolevel} 1000    5.0m 0.0  90.0)
*Vilo    2 0 sin(0.0 {lolevel} {rffreq} 5.0m 0.0  90.0)
Vilo     2 0 pulse(0.0 0.15 10.0m 2.0n 2.0n 71.43n 142.9n 0.0 )
Vqaudio 3 0 sin(0 {audiolevel} 1000    5.0m 0.0 0.0)
*Vqlo    4 0 sin(0.0 {lolevel} {rffreq} 5.0m 0.0 0.0)
Vqlo     4 0 pulse(0.0 0.15 10.0m 2.0n 2.0n 71.43n 142.9n 90.0 )


xampplusi  30 ampoutplusi  15 amplifier1
xampminusi 31 ampoutminusi 15 amplifier1

Lprimary1 ampoutplusi 15 500u
Lprimary2 15 ampoutminusi 500u
Lsecondary output 0 1000u
Ktrans1 Lprimary1 Lsecondary 1.0
Ktrans2 Lprimary2 Lsecondary 1.0
Ktrans3 Lprimary1 Lprimary2  1.0
Rload output 0 50.0

.control
set ngbehavior=ps

destroy all
save output ampoutplusi ampoutminusi 2 4

tran 2.0n 100.0m 90.0m uic

set lowlimit = 6.990e6
set highlimit = 7.010e6

plot v(ampoutplusi)
plot v(ampoutminusi)
plot v(2)
plot v(4)
plot v(output)

setplot tran1
linearize output
set specwindow = blackman 
fft output
plot db(output) xlimit $lowlimit $highlimit  ylimit -100 0.0 ydelta 10.0
plot db(output) ylimit -90.0 10.0 ydelta 10.0

.endc

.end
