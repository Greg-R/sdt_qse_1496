* Three Stage Power Amplifier Pre-Amplifier
* Include the sub-circuits.
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_original/simulation_first_stage/first_stage_amp_subckt.cir"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_original/simulation_second_stage/second_stage_amp_subckt.cir"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_original/simulation_third_stage/third_stage_subckt.cir"

* Power supply voltage source
Vsupply 15 0 15.0V

* Instantiate the 3 amplifier stages.
* Stage 1 has a resistive Pi attenuator on the input.  Blocking capacitor on output double normal value.
Xstage1 input output1 15  amplifier1
* Stage 2 has a blocking capacitor on the input which is double normal value.  No output blocking capacitor.
Xstage2     output1 output2 15  amplifier2
* Stage 3 has input and output blocking capacitors.
Xstage3 output2 output 15 amplifier3
*Rbig 2 0 1.0Meg
*Cout 2 output 0.1u


* Put a load on the output.
Rload output 0 100.0
Cload output 0 400p

.param audiolevel = 700m
*.param rffreq1 = 7.0Meg rffreq2 = 7.001Meg
.param rffreq1 = 7.0Meg rffreq2 = 7.001Meg

* Input signal source.
Vin1 10  0 sin(0 {audiolevel} {rffreq1} 10.0m 0 0)
* Another signal source in series for two-tone test.
Vin2 11  10 sin(0 {audiolevel} {rffreq2} 10.0m 0 0)
Rs  11 input 50.0

.control
set ngbehavior=ps
destroy all
save input output1 output2 output
*op
tran 4.0n 20.0m 10.0m

*plot v(input)
*plot v(output)
*plot v(output1)

setplot tran1
linearize output
set specwindow = blackman 
fft output
plot db(output) xlimit 6.995Meg 7.005Meg  ylimit -90 10.0 ydelta 10.0
*plot db(output) ylimit -90.0 10.0 ydelta 10.0

setplot tran1
linearize output1
set specwindow = blackman 
fft output1
plot db(output1) xlimit 6.995Meg 7.005Meg  ylimit -90 10.0 ydelta 10.0
*plot db(output1) ylimit -90.0 10.0 ydelta 10.0

setplot tran1
linearize output2
set specwindow = blackman 
fft output2
plot db(output2) xlimit 6.995Meg 7.005Meg  ylimit -90 10.0 ydelta 10.0
*plot db(output2) ylimit -90.0 10.0 ydelta 10.0

.endc

.end