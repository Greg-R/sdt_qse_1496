* Simulate MC1496 based IQ Modulator
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_iq_modulator/dsbmod_subckt.cir"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/feedback_amp_subckt.cir"

Vsupply 15 0 DC 12.27

* Modulator outputs are connected by thin transmission line.
xmodi 1 2 30 31 15 dsbmodulator
xmodq 3 4 30 31 15 dsbmodulator

* Add shunt capacitance to the modulator outputs.  This represents board stray capacitance.
Cmodstray1 30 0 0.001p
Comdstray2 31 0 0.001p

* DSB modulator output bias resistors
Rbiasi 15 30 510.0
Rbiasq 15 31 510.0

.param audiolevel = 100.0m lolevel = 150.0m
.param rffreq = 7.001e6

Viaudio 1 0 sin(0 {audiolevel} 1000    5.0m 0.0  90.0)
Vilo    2 0 sin(0.0 {lolevel} {rffreq} 5.0m 0.0  90.0)
*Vilo     2 0 pulse(0.0 0.05 150.0m 2.0n 2.0n 71.43n 142.9n 0.0 )
Vqaudio 3 0 sin(0 {audiolevel} 1000    5.0m 0.0 0.0)
Vqlo    4 0 sin(0.0 {lolevel} {rffreq} 5.0m 0.0 0.0)
*Vqlo     4 0 pulse(0.0 0.05 150.0m 2.0n 2.0n 71.43n 142.9n 90.0 )


*xampplusi  30 ampoutplusi  15 amplifier1
*xampminusi 31 ampoutminusi 15 amplifier1

* Output transformer
* Input leakage inductances
*Lleak1 ampoutplusi 32  0.03u
*Lleak2 ampoutminusi 33 0.03u
Lprimary1 30 15  32.0u
Lprimary2 15 31  32.0u
Lsecondary 34 0 32.0u
Lleakout 34 output     0.03u
Ktrans1 Lprimary1 Lsecondary 1.0
Ktrans2 Lprimary2 Lsecondary 1.0
Ktrans3 Lprimary1 Lprimary2  1.0
Rload output 0 50.0
*Cmatch output 0 75.0p

.control
set ngbehavior=ps

destroy all
save output ampoutplusi ampoutminusi v(30) v(31)

tran 2.0n 100.0m 90.0m uic

set lowlimit =  6.990e6
set highlimit = 7.010e6

plot v(ampoutplusi)
plot v(ampoutminusi)
plot v(30)
plot v(31)
plot v(output)

setplot tran1
linearize output
set specwindow = blackman 
fft output
plot db(output) xlimit $lowlimit $highlimit  ylimit -100 0.0 ydelta 10.0
plot db(output) ylimit -90.0 10.0 ydelta 10.0

.endc

.end
