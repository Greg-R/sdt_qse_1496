Simulate MC1496 based IQ Modulator
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/MC1496_SPICE_MODEL.LIB"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/MMBT2222ALT1.LIB"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_iq_modulator/dsbmod_subckt.cir"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/feedback_amp_subckt.cir"

xmodi 1 2 30 31 dsbmodulator
*xmodq 3 4 outplus outminus dsbmodulator

Vsupply 15 0 DC 12.27
*Qoutplusi  outplusQi 6 outplus Qmmbt2222alt1g
*Rplusload  15 outplusQi 100.0
*Rdiv1 15 6 1000.0
*Rdiv2  6 0 1000.0

.param audiolevel = 200.0m lolevel = 150.0m
.param rffreq = 28.0e6

Viaudio 1 0 sin(0 {audiolevel} 1000    5.0m 0.0  0)
Vilo    2 0 sin(0.0 {lolevel} {rffreq} 5.0m 0.0  0)
*Vqaudio 3 0 sin(0 {audiolevel} 1000    5.0m 0.0 90)
*Vqlo    4 0 sin(0.0 {lolevel} {rffreq} 5.0m 0.0 90)

* A transformer on the outout.
*CapI outplus 30 0.1u
*CapQ outminus 31 0.1u

xampi 30  ampoutplus  15 amplifier1
Rloadi ampoutplus 0 50.0
xampq 31 ampoutminus 15 amplifier1
Rloadq ampoutminus 0 50.0

*Lprimary 30 31 1000u
*Lsecondary output 0 25u
*Ktrans Lprimary Lsecondary 1.0

* RF Load
*Rload output 0 50.0

.control
set ngbehavior=ps

destroy all
save outplus outminus output ampoutplus ampoutminus

tran 2.0n 40.0m 30.0m uic
*setplot tran1
*plot output

set lowlimit = 27.995e6
set highlimit = 28.005e6

*let output  = (outplusi + outplusq) - (outminusi + outminusq)
*let output1 = outplusi - outminusi
*let output2 = outplusq - outminusq

*plot outplus
*plot outminus

plot v(ampoutplus)
plot v(ampoutminus)

let output = ampoutplus - ampoutminus
plot v(output)

*setplot tran1
*linearize output2
*set specwindow = blackman 
*fft output2
*plot db(output2) xlimit $lowlimit $highlimit  ylimit -90 10.0 ydelta 10.0
*plot db(output2) ylimit -90.0 10.0 ydelta 10.0

setplot tran1
linearize output
set specwindow = blackman 
fft output
plot db(output) xlimit $lowlimit $highlimit  ylimit -90 10.0 ydelta 10.0
plot db(output) ylimit -90.0 10.0 ydelta 10.0

*setplot tran1
*linearize xmodi.12
*set specwindow = blackman 
*fft xmodi.12
*plot db(xmodi.12) xlimit 6.995e6 7.005e6  ylimit -100 0.0 ydelta 10.0
*plot db(xmodi.12) ylimit -100.0 0.0 ydelta 10.0

.endc

.end
