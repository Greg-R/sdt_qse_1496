Simulate MC1496 based IQ Modulator
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation/MC1496_SPICE_MODEL.LIB"
.control
set ngbehavior=ps

save inaudio
save inrf
save output
save v(4)
save v(1)
save v(8)

tran 1n 20.1m
run

plot output
*plot v(8)
*plot v(4)
*plot v(1)
.endc

* MC1496 VS+ GAIN2 GAIN3 VS- Bias VO+ NC VEE NC VO- NC VC- NC VC+
XGCELL 1 2 3 4 5 6 7 0 9 12 11 10 13 8 MC1496

* 12 volt power supply

Vsupply 15 0 DC 12.27

* Output bias resistors
Rloadplus   15  6 3000
Rloadminus  15 12 3000

* Gain setting resistor
Rgain 2 3 1000

* Main bias control resistor
Rbias 15 5 10000

* Bias chain
R1 15  8 1300
R2  8 17  820
R3 17  0 1000

* Signal input bias
R4 17 1 1000
R5 17 4 1000

* Signal input blocking capacitor
C1 inaudio 1 0.1u

* Signal bypass capacitors, for both RF and audio.
Caudiobypass 4 0 100.0u
Crfbypass 8 0 100.0u

* Carrier input bias
R6 8 10 51

* Signal input and output blocking capacitors
C2 inrf 10 0.1u
Cout 6 output 0.01u
Rl output 0 10000

* Input excitation, 1 kHz tone.
Vaudio inaudio 0 sin(0 200m 1000 0.1m 0)

* Local Oscillator 7.0 MHz
Vlo inrf 0 Pulse(0.0, 0.0m, 0.1m, 2.0n, 2.0n, 7.1428e-8, 1.4286e-7)

.end
