*************************
      *from a web page
      *https://www.edaboard.com/threads/which-tool-can-simulate-mc1496.67325/
.subckt MC1496 1 2 3 4 5 6 8 10 12 14
* Tail current Source
Q1 3 5 19 Q2nn
Q2 2 5 13 Q2nn
* Input transistors
Q3 7 4 3 Q2nn
Q4 9 1 2 Q2nn
*LO quad switching Transistors
Q5 6 8 7 Q2nn
Q6 6 10 9 Q2nn
Q7 12 10 7 Q2nn
Q8 12 8 9 Q2nn
* Emitter degeneration resistors
RE1 19 14 500
RE2 13 14 500
*
* Current Mirror
Q9 5 5 15 Q2nn
Rd 15 14 500
.ENDS
.MODEL Q2nn NPN(
+ISS=0 XTF=1 NS=1
+CJS=0 VJS=0.5 PTF=0
+MJS=0 EG=1.1 AF=1
+ITF=0.5 VTF=1 BF=280.92203
+BR=20 IS=2.3673E-15 VAF=130.20848
+VAR=11.074004 IKF=0.23419 ISE=3.0707E-16
+NE=1.19409 IKR=7.80101 ISC=3.5223E-12
+NC=1.33867 IRB=1.8864E-4 NF=0.97302
+NR=0.97623 RBM=1E-2 RB=69.94226
+RC=3E-02 RE=0.2569 MJE=0.36064
+MJC=0.29228 VJE=0.81795 VJC=0.45460
+TF=5E-10 TR=6.2636E-09 CJE=6.7441E-12
+CJC=3.4247E-12 FC=0.95 XCJC=0.95425)
******************************************************
