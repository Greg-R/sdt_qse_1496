* Simulate a 2N3904 HF Amplifier
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_2N3904_amp/2N3904.LIB"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_xmas_travel/MMBT2222ALT1.LIB"

* Basic BJT biasing ...
*.options savecurrents

.subckt amplifier input output vsupply

*Q1 3 2 1 Q2n3904
Q1 3 2 1 Qmmbt2222alt1g

Rc  vsupply 5  100
Cc  5 0  0.1u
Lc  5 3  330u
R1  5 2  4700
R2  2 0  5100
R3  6 0   200
Rf  3 8   250
Cf  2 8  0.1u
Ci  input 2  0.1u
Re  1 6    10.0
Ce  6 0  0.1u
Co  3 output  0.1u

.ends amplifier