* Sub-circuit for the 1st Stage of the SDT Power Amplifier
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/2N3904.LIB"
*.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/MMBT2222ALT1.LIB"

* Basic BJT biasing ...
*.options savecurrents

.subckt amplifier1 input output vsupply

* NPN BJT Collector Base Emitter
Q1 vsupply 2 1 Q2n3904
*Q1 3 2 1 Qmmbt2222alt1g

* Input Pi attenuator.
R4 input 0   150.0
R17 input 12  37.0
R16 12  0 150.0

C1  12 2  0.1u

R1  vsupply 2  4700
R2  2 0        5100
R3  1 0         200

* Note that this coupling capacitor has double the capacitance.
* This is so when in series with the capacitor of the next stage the value will be correct.
C2 1 output 0.2u
Rbig output 0 2.0Meg

.ends amplifier1