* 2N3904 50 Ohm Amplifier Transient Test Bench

* Include the sub-circuit.
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_2N3904_amp/amplifier_2n3904.cir"

.param audiolevel = 400m
.param rffreq = 1.0Meg

* Instantiate an amplifier.
Xamplifier 1 2 3 amplifier

* Needs a 15 volt power source:
Vsupply 3 0 15V

Rload 2 0 50.0

* Input source
Vin 1 0 sin(0 {audiolevel} {rffreq} 0.1m 0 0)

.control
set ngbehavior=ps

*op
tran 20.0n 2.0m 1.99m

plot v(2)

.endc

.end

