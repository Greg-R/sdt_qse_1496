* Simulate a 2N3904 HF Amplifier
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/2N3904.LIB"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/MMBT2222ALT1.LIB"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/2sc4618.lib"

.subckt amplifier1 input output vsupply

*Q1 3 2 1 Q2n3904
*Q1 3 2 1 Qmmbt2222alt1g
Q1 output 2 1 Q2SC4618

*Rc  vsupply 5  100
*Cc  5 0  0.1u
*Lc  5 3  1000u
R1  vsupply 2  4700
R2  2 0  5100
R3  6 0   200
Rf  output 8   500
Cf  2 8  0.1u
Ci  input 2  0.1u
Re  1 6    10.0
Ce  6 0  0.1u
*Co  3 output  0.1u

*Rbig output 0 1Meg

.ends amplifier