Simulate MC1496 based IQ Modulator
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation/MC1496_SPICE_MODEL.LIB"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation/MMBT2222ALT1.LIB"

* 12 volt power supply
Vsupply 15 0 DC 12.27

.param audiolevel = 200m
.param lolevel    =  100m
.param rfload = 1000
.param remitter = 1000

* This is the I channel.
* MC1496 VS+ GAIN2 GAIN3 VS- Bias VO+ NC VEE NC VO- NC VC- NC VC+
XGCELL1 1 2 3 4 5 6 7 0 9 12 11 10 13 8 MC1496


* Begin 1st DSB modulator
* Output bias resistors
Rloadplusi   15  6 3000
Rloadminusi  15 12 3000
* Gain setting resistor
Rgain 2 3 1000
* Main bias control resistor
Rbias 15 5 10000
* Bias chain
R1 15  8 1300
R2  8 17  820
R3 17  0 1000
* Signal input bias
R4 17 1 1000
R5 17 4 1000
* Signal input blocking capacitor
C1i inaudio 1 0.1u
* Signal bypass capacitors, for both RF and audio.
Caudiobypassi 4 0 25.0u
Crfbypassi 8 0 25.0u
* Carrier input bias
R6i 8 10 51
* Signal input and output blocking capacitors
C2i inrf 10 0.1u
*Coutplusi 6 outputplusi 0.01u
*Rlplusi outputplusi 0 10000
*Coutminusi 12 outputminusi 0.01u
*Rlminusi outputminusi 0 10000

* Output emitter followers and blocking caps.
Qoutplusi  15 6 120 Qmmbt2222alt1g
Qoutminusi 15 12 121 Qmmbt2222alt1g
Rlplusi 120 0  remitter
Rlminusi 121 0 remitter
Coutplusi 120 outputplusi 0.1u
Coutminusi 121 outputminusi 0.1u

* Input excitation, 1 kHz tone.
Viaudio inaudio 0 sin(0 audiolevel 1000 0.1m 0 0)
* Local Oscillator 7.0 MHz
*Vilo inrf 0 Pulse(0.0, 50.0m, 0.1m, 2.0n, 2.0n, 0.5e-6, 1.0e-6)
Vilo inrf 0 sin(0.0, lolevel, 1.0e6, 0.1m, 0, 0)

* Begin 2nd DSB modulator which is the Q channel.
XGCELL2 101 102 103 104 105 106 107 0 109 112 111 110 113 108 MC1496
* Output bias resistors
Rloadplusq   15  106 3000
Rloadminusq  15 112 3000
* Gain setting resistor
Rgainq 102 103 1000
* Main bias control resistor
Rbiasq 15 105 10000
* Bias chain
R1q 15  108 1300
R2q  108 117  820
R3q 117  0 1000
* Signal input bias
R4q 117 101 1000
R5q 117 104 1000
* Signal input blocking capacitor
C1q qnaudio 101 0.1u
* Signal bypass capacitors, for both RF and audio.
Caudiobypassq 104 0 25.0u
Crfbypassq 108 0 25.0u
* Carrier input bias
R6q 108 110 51
* Signal input and output blocking capacitors
C2q qnrf 110 0.1u
*Coutplusq 112 outputplusq 0.01u
*Rlplusq   outputplusq 0 10000
*Coutminusq 106 outputminusq 0.01u
*Rlminusq outputminusq 0 10000

* Input excitation, 1 kHz tone.
Vqaudio qnaudio 0 sin(0 audiolevel 1000 0.1m 0 90)
* Local Oscillator 7.0 MHz
Vqlo qnrf 0 sin(0.0, lolevel, 1.0e6, 0.1m, 0 90)
*Vqlo qnrf 0 Pulse(0.0, 50.0m, 0.1m, 2.0n, 2.0n, 0.5e-6, 1.0e-6, 90)

* Output emitter followers and blocking capacitors.
Qoutplusq  15 106 122 Qmmbt2222alt1g
Qoutminusq 15 112 123 Qmmbt2222alt1g
Rlplusq 122 0  remitter
Rlminusq 123 0 remitter
Coutplusq 122 outputplusq 0.1u
Coutmniusq 123 outputminusq 0.1u

* Join the positive outputs together with small resistors.
Rplusi outputplusi outputplus 10
Rplusq outputplusq outputplus 10
Rloadplus outputplus 0 rfload

* Join the negative outputs together with small resistors.
Rminusi outputminusi outputminus 10
Rminusq outputminusq outputminus 10
Rloadminus outputminus 0 rfload

.control
*set ngbehavior=ps

destroy all
*set output = outputplus - outputminus
*save output twelve outputb



tran 20.0n 5.1m
*run

*plot outputi
*plot outputq
* v(6)
*plot v(106)
*plot output
*setplot tran1
*linearize output
*set specwindow = hamming
*fft output
*plot db(output) xlimit 0.995e6 1.005e6 ylimit -100 0.0 ydelta 10.0
*plot db(output) xlimit 0.0 20.0e6 ylimit -100 0.0 ydelta 10.0
*setplot tran1
*linearize twelve
*fft twelve
*plot db(twelve) xlimit 0.995e6 1.005e6 ylimit -100 0.0 ydelta 10.0
*let output = v(122) - v(123)
let output = outputplus - outputminus

plot output
*setplot tran1
*linearize output
*set specwindow = hamming
*fft output
*plot db(output) xlimit 0.995e6 1.005e6 ylimit -100 0.0 ydelta 10.0

*plot db(fft(output)) xlimit 0.995e6 1.005e6 ylimit -100 0.0 ydelta 10.0

*set bullshit = twelve
*set specwindow = blackman
*fft inaudio
*settype inaudio
*plot db(inaudio)

*plot inaudio qnaudio
*plot qnaudio
*plot inrf qnrf
*plot qnrf
*reset
.endc

.end
