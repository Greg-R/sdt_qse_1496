* 2N3904 50 Ohm Amplifier Test Bench

* Include the sub-circuit.
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_2N3904_amp/amplifier_2n3904.cir"

* Instantiate an amplifier.
Xamplifier 1 2 3 amplifier

* Needs a 15 volt power source:
Vsupply 3 0 15V

* Input source
Vin 1 0 dc 0 ac 1.0 portnum 1 z0 50.0
* Output source
Vout 2 0 dc 0 ac 1.0 portnum 2 z0 50.0


.control
set ngbehavior=ps
*op
*ac dec 10 1.0Meg 100.0Meg
sp dec 10 1.0Meg 100.0Meg

*plot vdb(7) xlog

.endc

.end

