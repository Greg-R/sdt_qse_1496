* Test of pulse transmformers.

Vsource 1 0 AC 1.0
Rsource 1 2 50.0

* Transformer
Linput 2 0 10.0u
Loutput 3 0 10.0u
Ktrans Linput Loutput 0.999

Rload 3 0 50.0


.control
save v(3)

ac dec 10 1.0Meg 30.0Meg

plot v(3)

.endc
.end