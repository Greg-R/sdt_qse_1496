* Simulate MC1496 based IQ Modulator.  Check the output impedance.
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/simulation_iq_modulator/dsbmod_subckt.cir"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/feedback_amp_subckt.cir"

Vsupply 15 0 DC 12.27

* Modulator outputs are connected by thin transmission line.
xmodi 1 2 30 31 15 dsbmodulator
xmodq 3 4 30 31 15 dsbmodulator

* Add shunt capacitance to the modulator outputs.  This represents board stray capacitance.
Cmodstray1 30 0 0.001p
Comdstray2 31 0 0.001p

* DSB modulator output bias resistors
Rbiasi 15 30 510.0
Rbiasq 15 31 510.0

*.param audiolevel = 100.0m lolevel = 150.0m
*.param rffreq = 28.001e6

* Put resistors in place of transient sources.
Riaduio 1 0 600.0
Rqaudio 3 0 600.0
Rilo    2 0 470.0
Rqlo    4 0 470.0

*Viaudio 1 0 sin(0 {audiolevel} 1000    5.0m 0.0  90.0)
*Vilo    2 0 sin(0.0 {lolevel} {rffreq} 5.0m 0.0  90.0)
*Vilo     2 0 pulse(0.0 0.05 150.0m 2.0n 2.0n 71.43n 142.9n 0.0 )
*Vqaudio 3 0 sin(0 {audiolevel} 1000    5.0m 0.0 0.0)
*Vqlo    4 0 sin(0.0 {lolevel} {rffreq} 5.0m 0.0 0.0)
*Vqlo     4 0 pulse(0.0 0.05 150.0m 2.0n 2.0n 71.43n 142.9n 90.0 )


xampplusi  30 ampoutplusi  15 amplifier1
xampminusi 31 ampoutminusi 15 amplifier1

* Output transformer
* Input leakage inductances
Lleak1 ampoutplusi 32  0.00003u
Lleak2 ampoutminusi 33 0.00003u
Lprimary1 32 15  32.0u
Lprimary2 15 33  32.0u
Lsecondary 34 0 32.0u
*Lleakout 34 output     0.00003u
Ktrans1 Lprimary1 Lsecondary 1.0
Ktrans2 Lprimary2 Lsecondary 1.0
Ktrans3 Lprimary1 Lprimary2  1.0
*Rload output 0 50.0
Cshunt 34 0 75.0p
*Lstry output 36 0.0005u
Vs22 34 0 portnum 2 z0 50.0

* Dummy port for Port 1
Rdummy 40 0 50.0
Ldummy 40 41 80.0n
Vs11   41 0 portnum 1 z0 50.0

.control
set ngbehavior=ps

destroy all
sp dec 10 3.0MEG 50.0MEG


plot s_2_2 smithgrid

*plot db(output) xlimit $lowlimit $highlimit  ylimit -100 0.0 ydelta 10.0
*plot db(output) ylimit -90.0 10.0 ydelta 10.0

.endc

.end
