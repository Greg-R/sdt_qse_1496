* Simulate a 2N3904 HF Amplifier
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/2N3904.LIB"
.include "/home/raven/gitrepos/pcb/sdt_qse_1496/model/MMBT2222ALT1.LIB"

* Basic BJT biasing ...
*.options savecurrents

.subckt amplifier1 input output vsupply

*Q1 3 2 1 Q2n3904
Q1 3 2 1 Qmmbt2222alt1g

* Input Pi attenuator.
*R4 input 0   150.0
*R17 input 12  37.0
*R16 12  0 150.0

Rc  vsupply 5  1
Cc  5 0  0.1u
Lc  5 3  1000u
R1  5 2  4700
R2  2 0  5100
R3  6 0   200
Rf  3 8   250
Cf  2 8  0.1u
Ci  input 2  0.1u
Re  1 6    10.0
Ce  6 0  0.1u
Co  3 output  0.2u

Rbig output 0 1Meg

.ends amplifier